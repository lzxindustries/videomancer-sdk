-- Videomancer SDK - Open source FPGA-based video effects development kit
-- Copyright (C) 2025 LZX Industries LLC
-- File: video_timing_pkg.vhd - Video Timing Package
-- License: GNU General Public License v3.0
-- https://github.com/lzxindustries/videomancer-sdk
--
-- This file is free software: you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
--
-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with this program. If not, see <https://www.gnu.org/licenses/>.
--
-- Description:
--   Constant data and types for video timing configurations.

--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package video_timing_pkg is

  constant C_VIDEO_TIMING_ID_WIDTH          : integer := 4;
  constant C_VIDEO_TIMING_ID_COUNT          : integer := (2 ** C_VIDEO_TIMING_ID_WIDTH);
  constant C_VIDEO_TIMING_DATA_WIDTH        : integer := 12;
  constant C_VIDEO_TIMING_ACCUMULATOR_WIDTH : integer := 16;

  subtype t_video_timing_id is std_logic_vector(C_VIDEO_TIMING_ID_WIDTH - 1 downto 0);

  constant C_NTSC      : t_video_timing_id := "0000"; -- 0
  constant C_PAL       : t_video_timing_id := "1000"; -- 8
  constant C_480P      : t_video_timing_id := "0100"; -- 4
  constant C_576P      : t_video_timing_id := "1100"; -- 12
  constant C_720P60    : t_video_timing_id := "1110"; -- 14
  constant C_720P5994  : t_video_timing_id := "0110"; -- 6
  constant C_720P50    : t_video_timing_id := "0101"; -- 5
  constant C_1080I60   : t_video_timing_id := "1010"; -- 10
  constant C_1080I5994 : t_video_timing_id := "0010"; -- 2
  constant C_1080I50   : t_video_timing_id := "0001"; -- 1
  constant C_1080P30   : t_video_timing_id := "0111"; -- 7
  constant C_1080P2997 : t_video_timing_id := "1101"; -- 13
  constant C_1080P25   : t_video_timing_id := "1011"; -- 11
  constant C_1080P24   : t_video_timing_id := "0011"; -- 3
  constant C_1080P2398 : t_video_timing_id := "1001"; -- 9

  type t_video_timing_port is record
    avid          : std_logic;
    hsync_n       : std_logic;
    vsync_n       : std_logic;
    field_n       : std_logic;
    vavid         : std_logic;
    hsync_start   : std_logic;
    vsync_start   : std_logic;
    avid_start    : std_logic;
    avid_end      : std_logic;
    is_interlaced : std_logic;
  end record;

  type t_video_stream_yuv444 is record
    y       : std_logic_vector(9 downto 0);
    u       : std_logic_vector(9 downto 0);
    v       : std_logic_vector(9 downto 0);
    avid    : std_logic;
    hsync_n : std_logic;
    vsync_n : std_logic;
    field_n : std_logic;
  end record;

  type t_video_stream_yuv422 is record
    y       : std_logic_vector(9 downto 0);
    c       : std_logic_vector(9 downto 0);
    avid    : std_logic;
    hsync_n : std_logic;
    vsync_n : std_logic;
    field_n : std_logic;
  end record;

  subtype t_video_timing_range is std_logic_vector(1 downto 0);

  constant C_ANIMATION  : t_video_timing_range := "00";
  constant C_VERTICAL   : t_video_timing_range := "01";
  constant C_HORIZONTAL : t_video_timing_range := "10";

  type t_video_timing_config is record
    clocks_per_line          : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    lines_per_frame          : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    frame_width              : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    frame_height             : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    -- -- havid_clks_1             : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    -- -- havid_clks_0             : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    -- -- vavid_a_clks_1           : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    -- -- vavid_a_lines_1          : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    -- -- vavid_a_clks_0           : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    -- -- vavid_a_lines_0          : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    -- -- vavid_b_clks_1           : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    -- -- vavid_b_lines_1          : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    -- -- vavid_b_clks_0           : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    -- -- vavid_b_lines_0          : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    -- -- field_clks_1             : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    -- -- field_lines_1            : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    -- -- field_clks_0             : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    -- -- field_lines_0            : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    fsync_clks               : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    fsync_lines              : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    hsync_clks_0             : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    hsync_clks_1             : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    hsync_clks_b_0           : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    hsync_clks_b_1           : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    csync_clks_0             : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    csync_clks_1             : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    csync_2x_a_clks_1        : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    csync_2x_a_clks_0        : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    csync_2x_b_clks_1        : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    csync_2x_b_clks_0        : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    eq_pulses_a_clks_1       : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    eq_pulses_a_lines_1      : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    eq_pulses_a_clks_0       : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    eq_pulses_a_lines_0      : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    eq_pulses_b_clks_1       : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    eq_pulses_b_lines_1      : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    eq_pulses_b_clks_0       : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    eq_pulses_b_lines_0      : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    csync_serration_a_clks_1 : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    csync_serration_a_clks_0 : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    csync_serration_b_clks_1 : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    csync_serration_b_clks_0 : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    csync_serration_c_clks_1 : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    csync_serration_c_clks_0 : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    csync_serration_d_clks_1 : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    csync_serration_d_clks_0 : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    vsync_a_clks_1           : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    vsync_a_lines_1          : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    vsync_a_clks_0           : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    vsync_a_lines_0          : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    vsync_b_clks_1           : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    vsync_b_lines_1          : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    vsync_b_clks_0           : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    vsync_b_lines_0          : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    trisync_en               : std_logic;
    hramp_increment          : unsigned(C_VIDEO_TIMING_ACCUMULATOR_WIDTH - 1 downto 0);
    vramp_increment          : unsigned(C_VIDEO_TIMING_ACCUMULATOR_WIDTH - 1 downto 0);
    top_field_first          : std_logic;
    is_interlaced            : std_logic;
    -- -- hsync_offset_hdmi_to_hdmi        : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    -- -- hsync_offset_hdmi_to_encoder     : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    -- -- hsync_offset_composite_to_hdmi        : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    -- -- hsync_offset_composite_to_encoder     : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    -- -- hsync_offset_component_to_hdmi        : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    -- -- hsync_offset_component_to_encoder     : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
    -- -- hsync_pulse_width        : unsigned(C_VIDEO_TIMING_DATA_WIDTH - 1 downto 0);
  end record;

  type t_video_timing_config_array is array (0 to C_VIDEO_TIMING_ID_COUNT - 1) of t_video_timing_config;

  constant C_VIDEO_TIMING_CONFIG_ARRAY : t_video_timing_config_array := (
    0                        => -- C_NTSC
    (clocks_per_line         => to_unsigned(858, C_VIDEO_TIMING_DATA_WIDTH),
    lines_per_frame          => to_unsigned(525, C_VIDEO_TIMING_DATA_WIDTH),
    frame_width              => to_unsigned(720, C_VIDEO_TIMING_DATA_WIDTH),
    frame_height             => to_unsigned(486, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_1            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_0            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_clks               => to_unsigned(858-38, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_lines              => to_unsigned(3, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_1             => to_unsigned(1 + 63, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_0             => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_1             => to_unsigned(1 + 63, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_0             => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_1        => to_unsigned(1 + 31, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_0        => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_1        => to_unsigned(1 + 429 + 31, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_0        => to_unsigned(1 + 429, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_0       => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_0      => to_unsigned(10, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_1       => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_1      => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_0       => to_unsigned(1 + 429, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_0      => to_unsigned(272, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_1       => to_unsigned(1 + 429, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_1      => to_unsigned(263, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_1 => to_unsigned(1 + 429 - 63, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_0 => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_1 => to_unsigned(1 + 858 - 63, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_0 => to_unsigned(1 + 429, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_1 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_0 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_1 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_0 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_0           => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_0          => to_unsigned(7, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_1           => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_1          => to_unsigned(4, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_0           => to_unsigned(1 + 429, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_0          => to_unsigned(269, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_1           => to_unsigned(1 + 429, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_1          => to_unsigned(266, C_VIDEO_TIMING_DATA_WIDTH),
    trisync_en               => '0',
    hramp_increment          => to_unsigned((2 ** C_VIDEO_TIMING_ACCUMULATOR_WIDTH) / 720, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    vramp_increment          => to_unsigned((2 ** C_VIDEO_TIMING_ACCUMULATOR_WIDTH) / 486, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    top_field_first          => '0',
    is_interlaced            => '1'
    -- hsync_offset_hdmi_to_hdmi        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_hdmi_to_encoder     => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_hdmi        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_encoder     => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_hdmi        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_encoder     => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_pulse_width        => to_unsigned(63, C_VIDEO_TIMING_DATA_WIDTH)
    ),
    8                        => -- C_PAL
    (clocks_per_line         => to_unsigned(864, C_VIDEO_TIMING_DATA_WIDTH),
    lines_per_frame          => to_unsigned(625, C_VIDEO_TIMING_DATA_WIDTH),
    frame_width              => to_unsigned(720, C_VIDEO_TIMING_DATA_WIDTH),
    frame_height             => to_unsigned(576, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_1            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_0            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_clks               => to_unsigned(864 - 38, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_lines              => to_unsigned(625, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_1             => to_unsigned(1 + 63, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_0             => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_1             => to_unsigned(1 + 63, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_0             => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_1        => to_unsigned(1 + 31, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_0        => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_1        => to_unsigned(1 + 432 + 31, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_0        => to_unsigned(1 + 432, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_0       => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_0      => to_unsigned(6, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_1       => to_unsigned(1 + 432, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_1      => to_unsigned(623, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_0       => to_unsigned(1 + 432, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_0      => to_unsigned(318, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_1       => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_1      => to_unsigned(311, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_1 => to_unsigned(1 + 432 - 63, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_0 => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_1 => to_unsigned(1 + 864 - 63, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_0 => to_unsigned(1 + 432, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_1 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_0 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_1 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_0 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_0           => to_unsigned(1 + 432, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_0          => to_unsigned(3, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_1           => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_1          => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_0           => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_0          => to_unsigned(316, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_1           => to_unsigned(1 + 432, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_1          => to_unsigned(313, C_VIDEO_TIMING_DATA_WIDTH),
    trisync_en               => '0',
    hramp_increment          => to_unsigned((2 ** C_VIDEO_TIMING_ACCUMULATOR_WIDTH) / 720, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    vramp_increment          => to_unsigned((2 ** C_VIDEO_TIMING_ACCUMULATOR_WIDTH) / 576, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    top_field_first          => '1',
    is_interlaced            => '1'
    -- hsync_offset_hdmi_to_hdmi        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_hdmi_to_encoder     => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_hdmi        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_encoder     => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_hdmi        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_encoder     => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_pulse_width        => to_unsigned(63, C_VIDEO_TIMING_DATA_WIDTH)
    ),
    4                        => -- C_480P
    (clocks_per_line         => to_unsigned(858, C_VIDEO_TIMING_DATA_WIDTH),
    lines_per_frame          => to_unsigned(525, C_VIDEO_TIMING_DATA_WIDTH),
    frame_width              => to_unsigned(720, C_VIDEO_TIMING_DATA_WIDTH),
    frame_height             => to_unsigned(480, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_1            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_0            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_clks               => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_lines              => to_unsigned(1 + 12, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_1             => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_0             => to_unsigned(1 + 63, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_1             => to_unsigned(1 + 63, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_0             => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_1        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_0        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_1        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_0        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_0       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_0      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_1       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_1      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_0       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_0      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_1       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_1      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_1 => to_unsigned(1 + 858 - 63, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_0 => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_1 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_0 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_1 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_0 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_1 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_0 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_0           => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_0          => to_unsigned(1 + 12, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_1           => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_1          => to_unsigned(1 + 6, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    trisync_en               => '0',
    hramp_increment          => to_unsigned((2 ** C_VIDEO_TIMING_ACCUMULATOR_WIDTH) / 720, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    vramp_increment          => to_unsigned((2 ** C_VIDEO_TIMING_ACCUMULATOR_WIDTH) / 480, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    top_field_first          => '1',
    is_interlaced            => '0'
    -- hsync_offset_hdmi_to_hdmi        => to_unsigned(858, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_hdmi_to_encoder     => to_unsigned(858, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_hdmi        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_encoder     => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_hdmi        => to_unsigned(858, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_encoder     => to_unsigned(858, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_pulse_width        => to_unsigned(63, C_VIDEO_TIMING_DATA_WIDTH)
    ),
    12                       => -- C_576P
    (clocks_per_line         => to_unsigned(864, C_VIDEO_TIMING_DATA_WIDTH),
    lines_per_frame          => to_unsigned(625, C_VIDEO_TIMING_DATA_WIDTH),
    frame_width              => to_unsigned(720, C_VIDEO_TIMING_DATA_WIDTH),
    frame_height             => to_unsigned(576, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_1            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_0            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_clks               => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_lines              => to_unsigned(1 + 10, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_1             => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_0             => to_unsigned(1 + 63, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_1             => to_unsigned(1 + 63, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_0             => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_1        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_0        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_1        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_0        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_0       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_0      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_1       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_1      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_0       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_0      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_1       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_1      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_1 => to_unsigned(1 + 864 - 63, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_0 => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_1 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_0 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_1 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_0 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_1 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_0 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_0           => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_0          => to_unsigned(1 + 10, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_1           => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_1          => to_unsigned(1 + 5, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    trisync_en               => '0',
    hramp_increment          => to_unsigned((2 ** C_VIDEO_TIMING_ACCUMULATOR_WIDTH) / 720, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    vramp_increment          => to_unsigned((2 ** C_VIDEO_TIMING_ACCUMULATOR_WIDTH) / 576, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    top_field_first          => '1',
    is_interlaced            => '0'
    -- hsync_offset_hdmi_to_hdmi        => to_unsigned(864, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_hdmi_to_encoder     => to_unsigned(864, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_hdmi        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_encoder     => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_hdmi        => to_unsigned(864, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_encoder     => to_unsigned(864, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_pulse_width        => to_unsigned(63, C_VIDEO_TIMING_DATA_WIDTH)
    ),
    14                       => -- C_720P60
    (clocks_per_line         => to_unsigned(1650, C_VIDEO_TIMING_DATA_WIDTH),
    lines_per_frame          => to_unsigned(750, C_VIDEO_TIMING_DATA_WIDTH),
    frame_width              => to_unsigned(1280, C_VIDEO_TIMING_DATA_WIDTH),
    frame_height             => to_unsigned(720, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_1            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_0            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_clks               => to_unsigned(1 + 1650 - 40 - 4, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_lines              => to_unsigned(4, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_1             => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_0             => to_unsigned(1 + 40, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_1             => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_0             => to_unsigned(1 + 1650 - 40, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_1        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_0        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_1        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_0        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_0       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_0      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_1       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_1      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_0       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_0      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_1       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_1      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_1 => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_0 => to_unsigned(1 + 40 + 220, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_1 => to_unsigned(1 + 1650 - 110, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_0 => to_unsigned(1 + 1650 - 40, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_1 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_0 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_1 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_0 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_0           => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_0          => to_unsigned(6, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_1           => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_1          => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    trisync_en               => '1',
    hramp_increment          => to_unsigned((2 ** C_VIDEO_TIMING_ACCUMULATOR_WIDTH) / 1280, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    vramp_increment          => to_unsigned((2 ** C_VIDEO_TIMING_ACCUMULATOR_WIDTH) / 720, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    top_field_first          => '1',
    is_interlaced            => '0'
    -- hsync_offset_hdmi_to_hdmi        => to_unsigned(1648, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_hdmi_to_encoder     => to_unsigned(1599, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_hdmi        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_encoder     => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_hdmi        => to_unsigned(1648, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_encoder     => to_unsigned(1605, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_pulse_width        => to_unsigned(40, C_VIDEO_TIMING_DATA_WIDTH)
    ),
    6                        => -- C_720P5994
    (clocks_per_line         => to_unsigned(1650, C_VIDEO_TIMING_DATA_WIDTH),
    lines_per_frame          => to_unsigned(750, C_VIDEO_TIMING_DATA_WIDTH),
    frame_width              => to_unsigned(1280, C_VIDEO_TIMING_DATA_WIDTH),
    frame_height             => to_unsigned(720, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_1            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_0            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_clks               => to_unsigned(1 + 1650 - 40 - 4, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_lines              => to_unsigned(4, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_1             => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_0             => to_unsigned(1 + 40, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_1             => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_0             => to_unsigned(1 + 1650 - 40, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_1        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_0        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_1        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_0        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_0       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_0      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_1       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_1      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_0       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_0      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_1       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_1      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_1 => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_0 => to_unsigned(1 + 40 + 220, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_1 => to_unsigned(1 + 1650 - 110, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_0 => to_unsigned(1 + 1650 - 40, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_1 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_0 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_1 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_0 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_0           => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_0          => to_unsigned(6, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_1           => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_1          => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    trisync_en               => '1',
    hramp_increment          => to_unsigned((2 ** C_VIDEO_TIMING_ACCUMULATOR_WIDTH) / 1280, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    vramp_increment          => to_unsigned((2 ** C_VIDEO_TIMING_ACCUMULATOR_WIDTH) / 720, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    top_field_first          => '1',
    is_interlaced            => '0'
    -- hsync_offset_hdmi_to_hdmi        => to_unsigned(1648, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_hdmi_to_encoder     => to_unsigned(1599, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_hdmi        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_encoder     => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_hdmi        => to_unsigned(1648, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_encoder     => to_unsigned(1605, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_pulse_width        => to_unsigned(40, C_VIDEO_TIMING_DATA_WIDTH)
    ),
    5                        => -- C_720P50
    (clocks_per_line         => to_unsigned(1980, C_VIDEO_TIMING_DATA_WIDTH),
    lines_per_frame          => to_unsigned(750, C_VIDEO_TIMING_DATA_WIDTH),
    frame_width              => to_unsigned(1280, C_VIDEO_TIMING_DATA_WIDTH),
    frame_height             => to_unsigned(720, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_1            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_0            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_clks               => to_unsigned(1 + 1980 - 40 - 4, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_lines              => to_unsigned(4, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_1             => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_0             => to_unsigned(1 + 40, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_1             => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_0             => to_unsigned(1 + 1980 - 40, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_1        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_0        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_1        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_0        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_0       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_0      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_1       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_1      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_0       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_0      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_1       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_1      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_1 => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_0 => to_unsigned(1 + 40 + 220, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_1 => to_unsigned(1 + 1980 - 110 - 328, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_0 => to_unsigned(1 + 1980 - 40, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_1 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_0 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_1 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_0 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_0           => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_0          => to_unsigned(6, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_1           => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_1          => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    trisync_en               => '1',
    hramp_increment          => to_unsigned((2 ** C_VIDEO_TIMING_ACCUMULATOR_WIDTH) / 1280, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    vramp_increment          => to_unsigned((2 ** C_VIDEO_TIMING_ACCUMULATOR_WIDTH) / 720, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    top_field_first          => '1',
    is_interlaced            => '0'
    -- hsync_offset_hdmi_to_hdmi        => to_unsigned(1978, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_hdmi_to_encoder     => to_unsigned(1929, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_hdmi        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_encoder     => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_hdmi        => to_unsigned(1978, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_encoder     => to_unsigned(1929, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_pulse_width        => to_unsigned(40, C_VIDEO_TIMING_DATA_WIDTH)
    ),
    10                       => -- C_1080I60
    (clocks_per_line         => to_unsigned(2200, C_VIDEO_TIMING_DATA_WIDTH),
    lines_per_frame          => to_unsigned(1125, C_VIDEO_TIMING_DATA_WIDTH),
    frame_width              => to_unsigned(1920, C_VIDEO_TIMING_DATA_WIDTH),
    frame_height             => to_unsigned(1080, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_1            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_0            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_clks               => to_unsigned(1 + 2200 - 44 + 1, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_lines              => to_unsigned(1125, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_1             => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_0             => to_unsigned(1 + 44, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_1           => to_unsigned(1 + 1100, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_0           => to_unsigned(1 + 1100 + 44, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_1             => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_0             => to_unsigned(1 + 2200 - 44, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_1        => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_0        => to_unsigned(1 + 1100 - 44, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_1        => to_unsigned(1 + 1100, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_0        => to_unsigned(1 + 2200 - 44, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_0       => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_0      => to_unsigned(7, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_1       => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_1      => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_0       => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_0      => to_unsigned(569, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_1       => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_1      => to_unsigned(563, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_1 => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_0 => to_unsigned(1 + 44 + 88, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_1 => to_unsigned(1 + 1100 - 88, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_0 => to_unsigned(1 + 1100 - 44, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_1 => to_unsigned(1 + 1100, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_0 => to_unsigned(1 + 1100 + 44 + 88, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_1 => to_unsigned(1 + 2200 - 88 , C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_0 => to_unsigned(1 + 2200 - 44, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_0           => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_0          => to_unsigned(6, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_1           => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_1          => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_0           => to_unsigned(1 + 1100, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_0          => to_unsigned(568, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_1           => to_unsigned(1 + 1100, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_1          => to_unsigned(563, C_VIDEO_TIMING_DATA_WIDTH),
    trisync_en               => '1',
    hramp_increment          => to_unsigned((2 ** C_VIDEO_TIMING_ACCUMULATOR_WIDTH) / 1920, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    vramp_increment          => to_unsigned((2 ** C_VIDEO_TIMING_ACCUMULATOR_WIDTH) / 1080, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    top_field_first          => '1',
    is_interlaced            => '1'
    -- hsync_offset_hdmi_to_hdmi        => to_unsigned(2198, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_hdmi_to_encoder     => to_unsigned(2149, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_hdmi        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_encoder     => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_hdmi        => to_unsigned(2198, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_encoder     => to_unsigned(2149, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_pulse_width        => to_unsigned(44, C_VIDEO_TIMING_DATA_WIDTH)
    ),
    2                        => -- C_1080I5994
    (clocks_per_line         => to_unsigned(2200, C_VIDEO_TIMING_DATA_WIDTH),
    lines_per_frame          => to_unsigned(1125, C_VIDEO_TIMING_DATA_WIDTH),
    frame_width              => to_unsigned(1920, C_VIDEO_TIMING_DATA_WIDTH),
    frame_height             => to_unsigned(1080, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_1            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_0            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_clks               => to_unsigned(1 + 2200 - 44 + 1, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_lines              => to_unsigned(1125, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_1             => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_0             => to_unsigned(1 + 44, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_1           => to_unsigned(1 + 1100, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_0           => to_unsigned(1 + 1100 + 44, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_1             => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_0             => to_unsigned(1 + 2200 - 44, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_1        => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_0        => to_unsigned(1 + 1100 - 44, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_1        => to_unsigned(1 + 1100, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_0        => to_unsigned(1 + 2200 - 44, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_0       => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_0      => to_unsigned(7, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_1       => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_1      => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_0       => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_0      => to_unsigned(569, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_1       => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_1      => to_unsigned(563, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_1 => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_0 => to_unsigned(1 + 44 + 88, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_1 => to_unsigned(1 + 1100 - 88, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_0 => to_unsigned(1 + 1100 - 44, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_1 => to_unsigned(1 + 1100, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_0 => to_unsigned(1 + 1100 + 44 + 88, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_1 => to_unsigned(1 + 2200 - 88 , C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_0 => to_unsigned(1 + 2200 - 44, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_0           => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_0          => to_unsigned(6, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_1           => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_1          => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_0           => to_unsigned(1 + 1100, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_0          => to_unsigned(568, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_1           => to_unsigned(1 + 1100, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_1          => to_unsigned(563, C_VIDEO_TIMING_DATA_WIDTH),
    trisync_en               => '1',
    hramp_increment          => to_unsigned((2 ** C_VIDEO_TIMING_ACCUMULATOR_WIDTH) / 1920, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    vramp_increment          => to_unsigned((2 ** C_VIDEO_TIMING_ACCUMULATOR_WIDTH) / 1080, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    top_field_first          => '1',
    is_interlaced            => '1'
    -- hsync_offset_hdmi_to_hdmi        => to_unsigned(2198, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_hdmi_to_encoder     => to_unsigned(2149, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_hdmi        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_encoder     => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_hdmi        => to_unsigned(2198, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_encoder     => to_unsigned(2149, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_pulse_width        => to_unsigned(44, C_VIDEO_TIMING_DATA_WIDTH
    ),
    1                        => -- C_1080I50
    (clocks_per_line         => to_unsigned(2640, C_VIDEO_TIMING_DATA_WIDTH),
    lines_per_frame          => to_unsigned(1125, C_VIDEO_TIMING_DATA_WIDTH),
    frame_width              => to_unsigned(1920, C_VIDEO_TIMING_DATA_WIDTH),
    frame_height             => to_unsigned(1080, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_1            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_0            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_clks               => to_unsigned(2640 - 44, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_lines              => to_unsigned(1125, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_1             => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_0             => to_unsigned(1 + 44, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_1           => to_unsigned(1 + 1320, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_0           => to_unsigned(1 + 1320 + 44, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_1             => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_0             => to_unsigned(1 + 2640 - 44, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_1        => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_0        => to_unsigned(1 + 1320 - 44, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_1        => to_unsigned(1 + 1320, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_0        => to_unsigned(1 + 2640 - 44, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_0       => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_0      => to_unsigned(7, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_1       => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_1      => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_0       => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_0      => to_unsigned(569, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_1       => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_1      => to_unsigned(563, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_1 => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_0 => to_unsigned(1 + 44 + 88, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_1 => to_unsigned(1 + 1320 - 88 - 220, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_0 => to_unsigned(1 + 1320 - 44, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_1 => to_unsigned(1 + 1320, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_0 => to_unsigned(1 + 1320 + 44 + 88, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_1 => to_unsigned(1 + 2640 - 88 - 220, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_0 => to_unsigned(1 + 2640 - 44, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_0           => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_0          => to_unsigned(6, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_1           => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_1          => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_0           => to_unsigned(1 + 1320, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_0          => to_unsigned(568, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_1           => to_unsigned(1 + 1320, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_1          => to_unsigned(563, C_VIDEO_TIMING_DATA_WIDTH),
    trisync_en               => '1',
    hramp_increment          => to_unsigned((2 ** C_VIDEO_TIMING_ACCUMULATOR_WIDTH) / 1920, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    vramp_increment          => to_unsigned((2 ** C_VIDEO_TIMING_ACCUMULATOR_WIDTH) / 1080, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    top_field_first          => '1',
    is_interlaced            => '1'
    -- hsync_offset_hdmi_to_hdmi        => to_unsigned(2638, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_hdmi_to_encoder     => to_unsigned(2589, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_hdmi        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_encoder     => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_hdmi        => to_unsigned(2638, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_encoder     => to_unsigned(2589, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_pulse_width        => to_unsigned(44, C_VIDEO_TIMING_DATA_WIDTH)
    ),
    7                        => -- C_1080P30
    (clocks_per_line         => to_unsigned(2200, C_VIDEO_TIMING_DATA_WIDTH),
    lines_per_frame          => to_unsigned(1125, C_VIDEO_TIMING_DATA_WIDTH),
    frame_width              => to_unsigned(1920, C_VIDEO_TIMING_DATA_WIDTH),
    frame_height             => to_unsigned(1080, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_1            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_0            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_clks               => to_unsigned(1 + 2200 - 44 + 1, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_lines              => to_unsigned(4, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_1             => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_0             => to_unsigned(1 + 44, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_1             => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_0             => to_unsigned(1 + 2200 - 44, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_1        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_0        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_1        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_0        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_0       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_0      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_1       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_1      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_0       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_0      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_1       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_1      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_1 => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_0 => to_unsigned(1 + 44 + 88, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_1 => to_unsigned(1 + 2200 - 88 , C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_0 => to_unsigned(1 + 2200 - 44, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_1 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_0 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_1 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_0 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_0           => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_0          => to_unsigned(6, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_1           => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_1          => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    trisync_en               => '1',
    hramp_increment          => to_unsigned((2 ** C_VIDEO_TIMING_ACCUMULATOR_WIDTH) / 1920, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    vramp_increment          => to_unsigned((2 ** C_VIDEO_TIMING_ACCUMULATOR_WIDTH) / 1080, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    top_field_first          => '1',
    is_interlaced            => '0'
    -- hsync_offset_hdmi_to_hdmi        => to_unsigned(2198, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_hdmi_to_encoder     => to_unsigned(2149, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_hdmi        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_encoder     => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_hdmi        => to_unsigned(2198, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_encoder     => to_unsigned(2149, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_pulse_width        => to_unsigned(44, C_VIDEO_TIMING_DATA_WIDTH)
    ),
    13                       => -- C_1080P2997
    (clocks_per_line         => to_unsigned(2200, C_VIDEO_TIMING_DATA_WIDTH),
    lines_per_frame          => to_unsigned(1125, C_VIDEO_TIMING_DATA_WIDTH),
    frame_width              => to_unsigned(1920, C_VIDEO_TIMING_DATA_WIDTH),
    frame_height             => to_unsigned(1080, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_1            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_0            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_clks               => to_unsigned(1 + 2200 - 44 + 1, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_lines              => to_unsigned(4, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_1             => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_0             => to_unsigned(1 + 44, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_1             => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_0             => to_unsigned(1 + 2200 - 44, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_1        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_0        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_1        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_0        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_0       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_0      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_1       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_1      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_0       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_0      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_1       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_1      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_1 => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_0 => to_unsigned(1 + 44 + 88, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_1 => to_unsigned(1 + 2200 - 88 , C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_0 => to_unsigned(1 + 2200 - 44, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_1 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_0 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_1 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_0 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_0           => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_0          => to_unsigned(6, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_1           => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_1          => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    trisync_en               => '1',
    hramp_increment          => to_unsigned((2 ** C_VIDEO_TIMING_ACCUMULATOR_WIDTH) / 1920, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    vramp_increment          => to_unsigned((2 ** C_VIDEO_TIMING_ACCUMULATOR_WIDTH) / 1080, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    top_field_first          => '1',
    is_interlaced            => '0'
    -- hsync_offset_hdmi_to_hdmi        => to_unsigned(2198, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_hdmi_to_encoder     => to_unsigned(2149, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_hdmi        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_encoder     => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_hdmi        => to_unsigned(2198, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_encoder     => to_unsigned(2149, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_pulse_width        => to_unsigned(44, C_VIDEO_TIMING_DATA_WIDTH)
    ),
    11                       => -- C_1080P25
    (clocks_per_line         => to_unsigned(2640, C_VIDEO_TIMING_DATA_WIDTH),
    lines_per_frame          => to_unsigned(1125, C_VIDEO_TIMING_DATA_WIDTH),
    frame_width              => to_unsigned(1920, C_VIDEO_TIMING_DATA_WIDTH),
    frame_height             => to_unsigned(1080, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_1            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_0            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_clks               => to_unsigned(1 + 2640 - 44 + 1, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_lines              => to_unsigned(4, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_1             => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_0             => to_unsigned(1 + 44, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_1             => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_0             => to_unsigned(1 + 2640 - 44, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_1        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_0        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_1        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_0        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_0       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_0      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_1       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_1      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_0       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_0      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_1       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_1      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_1 => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_0 => to_unsigned(1 + 44 + 88, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_1 => to_unsigned(1 + 2640 - 88 - 438, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_0 => to_unsigned(1 + 2640 - 44, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_1 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_0 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_1 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_0 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_0           => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_0          => to_unsigned(6, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_1           => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_1          => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    trisync_en               => '1',
    hramp_increment          => to_unsigned((2 ** C_VIDEO_TIMING_ACCUMULATOR_WIDTH) / 1920, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    vramp_increment          => to_unsigned((2 ** C_VIDEO_TIMING_ACCUMULATOR_WIDTH) / 1080, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    top_field_first          => '1',
    is_interlaced            => '0'
    -- hsync_offset_hdmi_to_hdmi        => to_unsigned(2638, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_hdmi_to_encoder     => to_unsigned(2589, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_hdmi        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_encoder     => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_hdmi        => to_unsigned(2638, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_encoder     => to_unsigned(2589, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_pulse_width        => to_unsigned(44, C_VIDEO_TIMING_DATA_WIDTH)
    ),
    3                        => -- C_1080P24
    (clocks_per_line         => to_unsigned(2750, C_VIDEO_TIMING_DATA_WIDTH),
    lines_per_frame          => to_unsigned(1125, C_VIDEO_TIMING_DATA_WIDTH),
    frame_width              => to_unsigned(1920, C_VIDEO_TIMING_DATA_WIDTH),
    frame_height             => to_unsigned(1080, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_1            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_0            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_clks               => to_unsigned(1 + 2750 - 44 + 1, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_lines              => to_unsigned(4, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_1             => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_0             => to_unsigned(1 + 44, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_1             => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_0             => to_unsigned(1 + 2750 - 44, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_1        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_0        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_1        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_0        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_0       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_0      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_1       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_1      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_0       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_0      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_1       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_1      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_1 => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_0 => to_unsigned(1 + 44 + 88, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_1 => to_unsigned(1 + 2750 - 88 - 548, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_0 => to_unsigned(1 + 2750 - 44, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_1 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_0 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_1 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_0 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_0           => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_0          => to_unsigned(6, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_1           => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_1          => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    trisync_en               => '1',
    hramp_increment          => to_unsigned((2 ** C_VIDEO_TIMING_ACCUMULATOR_WIDTH) / 1920, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    vramp_increment          => to_unsigned((2 ** C_VIDEO_TIMING_ACCUMULATOR_WIDTH) / 1080, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    top_field_first          => '1',
    is_interlaced            => '0'
    -- hsync_offset_hdmi_to_hdmi        => to_unsigned(2748, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_hdmi_to_encoder     => to_unsigned(2699, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_hdmi        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_encoder     => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_hdmi        => to_unsigned(2748, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_encoder     => to_unsigned(2699, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_pulse_width        => to_unsigned(44, C_VIDEO_TIMING_DATA_WIDTH)
    ),
    9                        => -- C_1080P2398
    (clocks_per_line         => to_unsigned(2750, C_VIDEO_TIMING_DATA_WIDTH),
    lines_per_frame          => to_unsigned(1125, C_VIDEO_TIMING_DATA_WIDTH),
    frame_width              => to_unsigned(1920, C_VIDEO_TIMING_DATA_WIDTH),
    frame_height             => to_unsigned(1080, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_1            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_0            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_clks               => to_unsigned(1 + 2750 - 44 + 1, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_lines              => to_unsigned(4, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_1             => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_0             => to_unsigned(1 + 44, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_1             => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_0             => to_unsigned(1 + 2750 - 44, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_1        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_0        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_1        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_0        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_0       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_0      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_1       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_1      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_0       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_0      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_1       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_1      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_1 => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_0 => to_unsigned(1 + 44 + 88, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_1 => to_unsigned(1 + 2750 - 88 - 548, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_0 => to_unsigned(1 + 2750 - 44, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_1 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_0 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_1 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_0 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_0           => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_0          => to_unsigned(6, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_1           => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_1          => to_unsigned(1, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    trisync_en               => '1',
    hramp_increment          => to_unsigned((2 ** C_VIDEO_TIMING_ACCUMULATOR_WIDTH) / 1920, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    vramp_increment          => to_unsigned((2 ** C_VIDEO_TIMING_ACCUMULATOR_WIDTH) / 1080, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    top_field_first          => '1',
    is_interlaced            => '0'
    -- hsync_offset_hdmi_to_hdmi        => to_unsigned(2748, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_hdmi_to_encoder     => to_unsigned(2699, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_hdmi        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_encoder     => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_hdmi        => to_unsigned(2748, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_encoder     => to_unsigned(2699, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_pulse_width        => to_unsigned(44, C_VIDEO_TIMING_DATA_WIDTH)
    ),
    others                   =>
    (clocks_per_line         => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    lines_per_frame          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    frame_width              => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    frame_height             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- havid_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_a_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- vavid_b_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_1            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- field_lines_0            => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_clks               => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    fsync_lines              => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    hsync_clks_b_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_1             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_clks_0             => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_1        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_a_clks_0        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_1        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_2x_b_clks_0        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_0       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_0      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_clks_1       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_a_lines_1      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_0       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_0      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_clks_1       => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    eq_pulses_b_lines_1      => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_1 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_a_clks_0 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_1 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_b_clks_0 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_1 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_c_clks_0 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_1 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    csync_serration_d_clks_0 => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_a_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_0           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_0          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_clks_1           => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    vsync_b_lines_1          => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    trisync_en               => '0',
    hramp_increment          => to_unsigned(0, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    vramp_increment          => to_unsigned(0, C_VIDEO_TIMING_ACCUMULATOR_WIDTH),
    top_field_first          => '1',
    is_interlaced            => '0'
    -- hsync_offset_hdmi_to_hdmi        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_hdmi_to_encoder     => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_hdmi        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_composite_to_encoder     => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_hdmi        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_offset_component_to_encoder     => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH),
    -- hsync_pulse_width        => to_unsigned(0, C_VIDEO_TIMING_DATA_WIDTH)
    )
  );

end package;
